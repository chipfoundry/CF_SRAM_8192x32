VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CF_SRAM_8192x32
  CLASS BLOCK ;
  FOREIGN CF_SRAM_8192x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1450.000 BY 920.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 20.940 5.200 22.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.940 438.010 22.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.940 878.005 22.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 70.940 5.200 72.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 70.940 438.010 72.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 70.940 878.005 72.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 120.940 5.200 122.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 120.940 438.010 122.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 120.940 878.005 122.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 170.940 5.200 172.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 170.940 438.010 172.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 170.940 878.005 172.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 220.940 5.200 222.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 220.940 438.010 222.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 220.940 878.005 222.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 270.940 5.200 272.700 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 270.940 438.150 272.700 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 270.940 878.145 272.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 320.940 5.200 322.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 320.940 438.010 322.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 320.940 878.005 322.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 370.940 5.200 372.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 370.940 438.010 372.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 370.940 878.005 372.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 420.940 5.200 422.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 420.940 438.010 422.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 420.940 878.005 422.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 470.940 5.200 472.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 470.940 438.010 472.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 470.940 878.005 472.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 520.940 5.200 522.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 520.940 438.010 522.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 520.940 878.005 522.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 570.940 5.200 572.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 570.940 438.010 572.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 570.940 878.005 572.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 620.940 5.200 622.700 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 620.940 438.150 622.700 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 620.940 878.145 622.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 670.940 5.200 672.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 670.940 438.010 672.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 670.940 878.005 672.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 720.940 5.200 722.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 720.940 438.010 722.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 720.940 878.005 722.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 770.940 5.200 772.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 770.940 438.010 772.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 770.940 878.005 772.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 820.940 5.200 822.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 820.940 438.010 822.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 820.940 878.005 822.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 870.940 5.200 872.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 870.940 438.010 872.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 870.940 878.005 872.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 920.940 5.200 922.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 920.940 438.010 922.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 920.940 878.005 922.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 970.940 5.200 972.700 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 970.940 438.150 972.700 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 970.940 878.145 972.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1020.940 5.200 1022.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1020.940 438.010 1022.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1020.940 878.005 1022.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1070.940 5.200 1072.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1070.940 438.010 1072.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1070.940 878.005 1072.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1120.940 5.200 1122.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1120.940 438.010 1122.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1120.940 878.005 1122.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1170.940 5.200 1172.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1170.940 438.010 1172.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1170.940 878.005 1172.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1220.940 5.200 1222.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1220.940 438.010 1222.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1220.940 878.005 1222.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1270.940 5.200 1272.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1270.940 438.010 1272.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1270.940 878.005 1272.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1320.940 5.200 1322.700 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 1320.940 438.150 1322.700 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 1320.940 878.145 1322.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1370.940 5.200 1372.700 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1370.940 438.010 1372.700 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1370.940 878.005 1372.700 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1420.940 5.200 1422.700 914.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 21.320 1445.100 23.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 71.320 1445.100 73.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 121.320 1445.100 123.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 171.320 1445.100 173.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 221.320 1445.100 223.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 271.320 1445.100 273.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 321.320 1445.100 323.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 371.320 1445.100 373.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 421.320 1445.100 423.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 471.320 1445.100 473.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 521.320 1445.100 523.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 571.320 1445.100 573.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 621.320 1445.100 623.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 721.320 1445.100 723.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 771.320 1445.100 773.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 821.320 1445.100 823.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 871.320 1445.100 873.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.990 671.320 349.800 673.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 674.990 671.320 699.800 673.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1024.990 671.320 1049.800 673.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1374.990 671.320 1445.100 673.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.510 0.000 26.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.510 0.000 56.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.510 0.000 86.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.510 0.000 116.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.510 0.000 146.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.510 0.000 176.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.510 0.000 206.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.510 0.000 236.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.510 0.000 266.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.510 0.000 296.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.510 0.000 326.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 353.510 0.000 356.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.510 0.000 386.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.510 0.000 416.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.510 0.000 446.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.510 0.000 476.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.510 0.000 506.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.510 0.000 536.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.510 0.000 566.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.510 0.000 596.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.510 0.000 626.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.510 0.000 656.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.510 0.000 686.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 713.510 0.000 716.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.510 0.000 746.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.510 0.000 776.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.510 0.000 806.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 833.510 0.000 836.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.510 0.000 866.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 893.510 0.000 896.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.510 0.000 926.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.510 0.000 956.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 983.510 0.000 986.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.510 0.000 1016.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1043.510 0.000 1046.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.510 0.000 1076.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.510 0.000 1106.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1133.510 0.000 1136.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.510 0.000 1166.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1193.510 0.000 1196.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.510 0.000 1226.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1253.510 0.000 1256.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.510 0.000 1286.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1313.510 0.000 1316.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1343.510 0.000 1346.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.510 0.000 1376.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.510 0.000 1406.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1433.510 0.000 1436.610 920.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 331.930 26.960 333.690 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 681.530 464.880 683.290 881.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 331.930 464.880 333.690 881.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 681.530 26.960 683.290 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 1031.590 26.960 1033.350 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 1031.590 464.880 1033.350 881.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 453.020 1422.700 454.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 895.020 1422.700 896.780 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 9.180 5.200 10.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.180 438.150 10.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.180 878.145 10.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.180 5.200 60.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.180 438.010 60.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.180 878.005 60.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 109.180 5.200 110.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 109.180 438.010 110.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 109.180 878.005 110.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 159.180 5.200 160.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 159.180 438.010 160.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 159.180 878.005 160.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.180 5.200 210.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.180 438.010 210.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.180 878.005 210.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 259.180 5.200 260.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 259.180 438.150 260.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 259.180 878.145 260.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 309.180 5.200 310.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 309.180 438.010 310.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 309.180 878.005 310.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 359.180 5.200 360.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 359.180 438.150 360.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 359.180 878.145 360.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 409.180 5.200 410.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 409.180 438.010 410.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 409.180 878.005 410.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 459.180 5.200 460.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 459.180 438.010 460.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 459.180 878.005 460.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 509.180 5.200 510.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 509.180 438.010 510.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 509.180 878.005 510.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 559.180 5.200 560.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 559.180 438.010 560.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 559.180 878.005 560.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 609.180 5.200 610.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 609.180 438.150 610.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 609.180 878.145 610.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 659.180 5.200 660.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 659.180 438.010 660.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 659.180 878.005 660.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 709.180 5.200 710.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 709.180 438.150 710.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 709.180 878.145 710.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 759.180 5.200 760.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 759.180 438.010 760.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 759.180 878.005 760.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 809.180 5.200 810.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 809.180 438.010 810.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 809.180 878.005 810.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 859.180 5.200 860.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 859.180 438.010 860.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 859.180 878.005 860.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 909.180 5.200 910.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 909.180 438.010 910.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 909.180 878.005 910.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 959.180 5.200 960.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 959.180 438.150 960.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 959.180 878.145 960.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1009.180 5.200 1010.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1009.180 438.010 1010.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1009.180 878.005 1010.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1059.180 5.200 1060.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 1059.180 438.150 1060.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 1059.180 878.145 1060.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1109.180 5.200 1110.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1109.180 438.010 1110.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1109.180 878.005 1110.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1159.180 5.200 1160.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1159.180 438.010 1160.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1159.180 878.005 1160.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1209.180 5.200 1210.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1209.180 438.010 1210.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1209.180 878.005 1210.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1259.180 5.200 1260.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1259.180 438.010 1260.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1259.180 878.005 1260.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1309.180 5.200 1310.940 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 1309.180 438.150 1310.940 469.715 ;
    END
    PORT
      LAYER met2 ;
        RECT 1309.180 878.145 1310.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1359.180 5.200 1360.940 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1359.180 438.010 1360.940 469.855 ;
    END
    PORT
      LAYER met2 ;
        RECT 1359.180 878.005 1360.940 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 1409.180 5.200 1410.940 914.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 9.560 1445.100 11.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 59.560 1445.100 61.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 109.560 1445.100 111.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 159.560 1445.100 161.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 209.560 1445.100 211.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 259.560 1445.100 261.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 309.560 1445.100 311.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 359.560 1445.100 361.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 409.560 1445.100 411.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 459.560 1445.100 461.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 509.560 1445.100 511.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 559.560 1445.100 561.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 609.560 1445.100 611.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 659.560 1445.100 661.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 709.560 1445.100 711.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 759.560 1445.100 761.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 809.560 1445.100 811.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 859.560 1445.100 861.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.820 909.560 1445.100 911.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.510 0.000 11.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.510 0.000 41.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.510 0.000 71.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.510 0.000 101.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.510 0.000 131.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.510 0.000 161.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.510 0.000 191.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.510 0.000 221.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.510 0.000 251.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.510 0.000 281.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.510 0.000 311.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.510 0.000 341.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.510 0.000 371.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 398.510 0.000 401.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.510 0.000 431.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.510 0.000 461.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.510 0.000 491.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.510 0.000 521.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.510 0.000 551.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 578.510 0.000 581.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.510 0.000 611.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.510 0.000 641.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.510 0.000 671.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 698.510 0.000 701.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.510 0.000 731.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.510 0.000 761.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 788.510 0.000 791.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.510 0.000 821.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.510 0.000 851.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 878.510 0.000 881.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.510 0.000 911.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 938.510 0.000 941.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 968.510 0.000 971.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.510 0.000 1001.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1028.510 0.000 1031.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.510 0.000 1061.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.510 0.000 1091.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1118.510 0.000 1121.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1148.510 0.000 1151.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.510 0.000 1181.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.510 0.000 1211.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1238.510 0.000 1241.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.510 0.000 1271.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1298.510 0.000 1301.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1328.510 0.000 1331.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.510 0.000 1361.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1388.510 0.000 1391.610 920.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1418.510 0.000 1421.610 920.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 343.890 26.960 345.650 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 693.490 464.880 695.250 881.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 343.890 464.880 345.650 881.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 693.490 26.960 695.250 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 1043.550 26.960 1045.310 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 1043.550 464.880 1045.310 881.520 ;
    END
  END VPWR
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.150 0.000 971.430 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.130 0.000 1000.410 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 0.000 1116.330 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 0.000 1174.290 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.990 0.000 1203.270 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.970 0.000 1232.250 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.950 0.000 1261.230 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.930 0.000 1290.210 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.890 0.000 1348.170 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.870 0.000 1377.150 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 806.930 0.000 807.210 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 835.910 0.000 836.190 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 864.890 0.000 865.170 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 951.830 0.000 952.110 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1038.770 0.000 1039.050 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1067.750 0.000 1068.030 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1096.730 0.000 1097.010 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1154.690 0.000 1154.970 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1212.650 0.000 1212.930 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1241.630 0.000 1241.910 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1270.610 0.000 1270.890 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1328.570 0.000 1328.850 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1386.530 0.000 1386.810 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1415.510 0.000 1415.790 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 816.590 0.000 816.870 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 874.550 0.000 874.830 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 990.470 0.000 990.750 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1019.450 0.000 1019.730 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1106.390 0.000 1106.670 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1135.370 0.000 1135.650 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1193.330 0.000 1193.610 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1222.310 0.000 1222.590 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1251.290 0.000 1251.570 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1280.270 0.000 1280.550 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1309.250 0.000 1309.530 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1338.230 0.000 1338.510 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1367.210 0.000 1367.490 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 565.430 0.000 565.710 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1396.190 0.000 1396.470 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1425.170 0.000 1425.450 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 4.870 5.320 1445.050 914.005 ;
      LAYER li1 ;
        RECT 5.060 5.355 1444.860 914.005 ;
      LAYER met1 ;
        RECT 5.060 0.040 1444.860 914.160 ;
      LAYER met2 ;
        RECT 10.130 470.135 331.650 868.690 ;
        RECT 10.130 469.995 20.660 470.135 ;
        RECT 11.220 437.870 20.660 469.995 ;
        RECT 10.130 437.730 20.660 437.870 ;
        RECT 22.980 437.730 58.900 470.135 ;
        RECT 61.220 437.730 70.660 470.135 ;
        RECT 72.980 437.730 108.900 470.135 ;
        RECT 111.220 437.730 120.660 470.135 ;
        RECT 122.980 437.730 158.900 470.135 ;
        RECT 161.220 437.730 170.660 470.135 ;
        RECT 172.980 437.730 208.900 470.135 ;
        RECT 211.220 437.730 220.660 470.135 ;
        RECT 222.980 469.995 308.900 470.135 ;
        RECT 222.980 437.870 258.900 469.995 ;
        RECT 261.220 437.870 270.660 469.995 ;
        RECT 272.980 437.870 308.900 469.995 ;
        RECT 222.980 437.730 308.900 437.870 ;
        RECT 311.220 437.730 320.660 470.135 ;
        RECT 322.980 464.600 331.650 470.135 ;
        RECT 333.970 464.600 343.610 868.690 ;
        RECT 345.930 470.135 681.250 868.690 ;
        RECT 345.930 469.995 370.660 470.135 ;
        RECT 345.930 464.600 358.900 469.995 ;
        RECT 322.980 441.160 358.900 464.600 ;
        RECT 322.980 437.730 331.650 441.160 ;
        RECT 10.130 30.140 331.650 437.730 ;
        RECT 10.130 30.000 20.660 30.140 ;
        RECT 11.220 4.920 20.660 30.000 ;
        RECT 22.980 4.920 58.900 30.140 ;
        RECT 61.220 4.920 70.660 30.140 ;
        RECT 72.980 4.920 108.900 30.140 ;
        RECT 111.220 4.920 120.660 30.140 ;
        RECT 122.980 4.920 158.900 30.140 ;
        RECT 161.220 4.920 170.660 30.140 ;
        RECT 172.980 4.920 208.900 30.140 ;
        RECT 211.220 4.920 220.660 30.140 ;
        RECT 222.980 30.000 308.900 30.140 ;
        RECT 222.980 4.920 258.900 30.000 ;
        RECT 261.220 4.920 270.660 30.000 ;
        RECT 272.980 4.920 308.900 30.000 ;
        RECT 311.220 4.920 320.660 30.140 ;
        RECT 322.980 26.680 331.650 30.140 ;
        RECT 333.970 26.680 343.610 441.160 ;
        RECT 345.930 437.870 358.900 441.160 ;
        RECT 361.220 437.870 370.660 469.995 ;
        RECT 345.930 437.730 370.660 437.870 ;
        RECT 372.980 437.730 408.900 470.135 ;
        RECT 411.220 437.730 420.660 470.135 ;
        RECT 422.980 437.730 458.900 470.135 ;
        RECT 461.220 437.730 470.660 470.135 ;
        RECT 472.980 437.730 508.900 470.135 ;
        RECT 511.220 437.730 520.660 470.135 ;
        RECT 522.980 437.730 558.900 470.135 ;
        RECT 561.220 437.730 570.660 470.135 ;
        RECT 572.980 469.995 658.900 470.135 ;
        RECT 572.980 437.870 608.900 469.995 ;
        RECT 611.220 437.870 620.660 469.995 ;
        RECT 622.980 437.870 658.900 469.995 ;
        RECT 572.980 437.730 658.900 437.870 ;
        RECT 661.220 437.730 670.660 470.135 ;
        RECT 672.980 464.600 681.250 470.135 ;
        RECT 683.570 464.600 693.210 868.690 ;
        RECT 695.530 470.135 1031.310 868.690 ;
        RECT 695.530 469.995 720.660 470.135 ;
        RECT 695.530 464.600 708.900 469.995 ;
        RECT 672.980 441.160 708.900 464.600 ;
        RECT 672.980 437.730 681.250 441.160 ;
        RECT 345.930 30.140 681.250 437.730 ;
        RECT 345.930 30.000 370.660 30.140 ;
        RECT 345.930 26.680 358.900 30.000 ;
        RECT 322.980 4.920 358.900 26.680 ;
        RECT 361.220 4.920 370.660 30.000 ;
        RECT 372.980 4.920 408.900 30.140 ;
        RECT 411.220 4.920 420.660 30.140 ;
        RECT 422.980 4.920 458.900 30.140 ;
        RECT 461.220 4.920 470.660 30.140 ;
        RECT 472.980 4.920 508.900 30.140 ;
        RECT 511.220 4.920 520.660 30.140 ;
        RECT 522.980 4.920 558.900 30.140 ;
        RECT 561.220 4.920 570.660 30.140 ;
        RECT 572.980 30.000 658.900 30.140 ;
        RECT 572.980 4.920 608.900 30.000 ;
        RECT 611.220 4.920 620.660 30.000 ;
        RECT 622.980 4.920 658.900 30.000 ;
        RECT 661.220 4.920 670.660 30.140 ;
        RECT 672.980 26.680 681.250 30.140 ;
        RECT 683.570 26.680 693.210 441.160 ;
        RECT 695.530 437.870 708.900 441.160 ;
        RECT 711.220 437.870 720.660 469.995 ;
        RECT 695.530 437.730 720.660 437.870 ;
        RECT 722.980 437.730 758.900 470.135 ;
        RECT 761.220 437.730 770.660 470.135 ;
        RECT 772.980 437.730 808.900 470.135 ;
        RECT 811.220 437.730 820.660 470.135 ;
        RECT 822.980 437.730 858.900 470.135 ;
        RECT 861.220 437.730 870.660 470.135 ;
        RECT 872.980 437.730 908.900 470.135 ;
        RECT 911.220 437.730 920.660 470.135 ;
        RECT 922.980 469.995 1008.900 470.135 ;
        RECT 922.980 437.870 958.900 469.995 ;
        RECT 961.220 437.870 970.660 469.995 ;
        RECT 972.980 437.870 1008.900 469.995 ;
        RECT 922.980 437.730 1008.900 437.870 ;
        RECT 1011.220 437.730 1020.660 470.135 ;
        RECT 1022.980 464.600 1031.310 470.135 ;
        RECT 1033.630 464.600 1043.270 868.690 ;
        RECT 1045.590 470.135 1408.900 868.690 ;
        RECT 1045.590 469.995 1070.660 470.135 ;
        RECT 1045.590 464.600 1058.900 469.995 ;
        RECT 1022.980 441.160 1058.900 464.600 ;
        RECT 1022.980 437.730 1031.310 441.160 ;
        RECT 695.530 30.140 1031.310 437.730 ;
        RECT 695.530 30.000 720.660 30.140 ;
        RECT 695.530 26.680 708.900 30.000 ;
        RECT 672.980 4.920 708.900 26.680 ;
        RECT 711.220 4.920 720.660 30.000 ;
        RECT 722.980 4.920 758.900 30.140 ;
        RECT 761.220 4.920 770.660 30.140 ;
        RECT 772.980 4.920 808.900 30.140 ;
        RECT 811.220 4.920 820.660 30.140 ;
        RECT 822.980 4.920 858.900 30.140 ;
        RECT 861.220 4.920 870.660 30.140 ;
        RECT 872.980 4.920 908.900 30.140 ;
        RECT 911.220 4.920 920.660 30.140 ;
        RECT 922.980 30.000 1008.900 30.140 ;
        RECT 922.980 4.920 958.900 30.000 ;
        RECT 961.220 4.920 970.660 30.000 ;
        RECT 972.980 4.920 1008.900 30.000 ;
        RECT 1011.220 4.920 1020.660 30.140 ;
        RECT 1022.980 26.680 1031.310 30.140 ;
        RECT 1033.630 26.680 1043.270 441.160 ;
        RECT 1045.590 437.870 1058.900 441.160 ;
        RECT 1061.220 437.870 1070.660 469.995 ;
        RECT 1045.590 437.730 1070.660 437.870 ;
        RECT 1072.980 437.730 1108.900 470.135 ;
        RECT 1111.220 437.730 1120.660 470.135 ;
        RECT 1122.980 437.730 1158.900 470.135 ;
        RECT 1161.220 437.730 1170.660 470.135 ;
        RECT 1172.980 437.730 1208.900 470.135 ;
        RECT 1211.220 437.730 1220.660 470.135 ;
        RECT 1222.980 437.730 1258.900 470.135 ;
        RECT 1261.220 437.730 1270.660 470.135 ;
        RECT 1272.980 469.995 1358.900 470.135 ;
        RECT 1272.980 437.870 1308.900 469.995 ;
        RECT 1311.220 437.870 1320.660 469.995 ;
        RECT 1322.980 437.870 1358.900 469.995 ;
        RECT 1272.980 437.730 1358.900 437.870 ;
        RECT 1361.220 437.730 1370.660 470.135 ;
        RECT 1372.980 437.730 1408.900 470.135 ;
        RECT 1045.590 30.140 1408.900 437.730 ;
        RECT 1045.590 30.000 1070.660 30.140 ;
        RECT 1045.590 26.680 1058.900 30.000 ;
        RECT 1022.980 4.920 1058.900 26.680 ;
        RECT 1061.220 4.920 1070.660 30.000 ;
        RECT 1072.980 4.920 1108.900 30.140 ;
        RECT 1111.220 4.920 1120.660 30.140 ;
        RECT 1122.980 4.920 1158.900 30.140 ;
        RECT 1161.220 4.920 1170.660 30.140 ;
        RECT 1172.980 4.920 1208.900 30.140 ;
        RECT 1211.220 4.920 1220.660 30.140 ;
        RECT 1222.980 4.920 1258.900 30.140 ;
        RECT 1261.220 4.920 1270.660 30.140 ;
        RECT 1272.980 30.000 1358.900 30.140 ;
        RECT 1272.980 4.920 1308.900 30.000 ;
        RECT 1311.220 4.920 1320.660 30.000 ;
        RECT 1322.980 4.920 1358.900 30.000 ;
        RECT 1361.220 4.920 1370.660 30.140 ;
        RECT 1372.980 4.920 1408.900 30.140 ;
        RECT 1411.220 4.920 1420.660 868.690 ;
        RECT 1422.980 4.920 1425.440 868.690 ;
        RECT 10.130 4.280 1425.440 4.920 ;
        RECT 10.130 0.010 410.590 4.280 ;
        RECT 411.430 0.010 420.250 4.280 ;
        RECT 421.090 0.010 429.910 4.280 ;
        RECT 430.750 0.010 439.570 4.280 ;
        RECT 440.410 0.010 449.230 4.280 ;
        RECT 450.070 0.010 458.890 4.280 ;
        RECT 459.730 0.010 468.550 4.280 ;
        RECT 469.390 0.010 478.210 4.280 ;
        RECT 479.050 0.010 487.870 4.280 ;
        RECT 488.710 0.010 497.530 4.280 ;
        RECT 498.370 0.010 507.190 4.280 ;
        RECT 508.030 0.010 516.850 4.280 ;
        RECT 517.690 0.010 526.510 4.280 ;
        RECT 527.350 0.010 536.170 4.280 ;
        RECT 537.010 0.010 545.830 4.280 ;
        RECT 546.670 0.010 555.490 4.280 ;
        RECT 556.330 0.010 565.150 4.280 ;
        RECT 565.990 0.010 574.810 4.280 ;
        RECT 575.650 0.010 584.470 4.280 ;
        RECT 585.310 0.010 594.130 4.280 ;
        RECT 594.970 0.010 603.790 4.280 ;
        RECT 604.630 0.010 613.450 4.280 ;
        RECT 614.290 0.010 623.110 4.280 ;
        RECT 623.950 0.010 632.770 4.280 ;
        RECT 633.610 0.010 642.430 4.280 ;
        RECT 643.270 0.010 652.090 4.280 ;
        RECT 652.930 0.010 661.750 4.280 ;
        RECT 662.590 0.010 671.410 4.280 ;
        RECT 672.250 0.010 681.070 4.280 ;
        RECT 681.910 0.010 690.730 4.280 ;
        RECT 691.570 0.010 700.390 4.280 ;
        RECT 701.230 0.010 710.050 4.280 ;
        RECT 710.890 0.010 719.710 4.280 ;
        RECT 720.550 0.010 729.370 4.280 ;
        RECT 730.210 0.010 739.030 4.280 ;
        RECT 739.870 0.010 748.690 4.280 ;
        RECT 749.530 0.010 758.350 4.280 ;
        RECT 759.190 0.010 768.010 4.280 ;
        RECT 768.850 0.010 777.670 4.280 ;
        RECT 778.510 0.010 787.330 4.280 ;
        RECT 788.170 0.010 796.990 4.280 ;
        RECT 797.830 0.010 806.650 4.280 ;
        RECT 807.490 0.010 816.310 4.280 ;
        RECT 817.150 0.010 825.970 4.280 ;
        RECT 826.810 0.010 835.630 4.280 ;
        RECT 836.470 0.010 845.290 4.280 ;
        RECT 846.130 0.010 854.950 4.280 ;
        RECT 855.790 0.010 864.610 4.280 ;
        RECT 865.450 0.010 874.270 4.280 ;
        RECT 875.110 0.010 883.930 4.280 ;
        RECT 884.770 0.010 893.590 4.280 ;
        RECT 894.430 0.010 903.250 4.280 ;
        RECT 904.090 0.010 912.910 4.280 ;
        RECT 913.750 0.010 922.570 4.280 ;
        RECT 923.410 0.010 932.230 4.280 ;
        RECT 933.070 0.010 941.890 4.280 ;
        RECT 942.730 0.010 951.550 4.280 ;
        RECT 952.390 0.010 961.210 4.280 ;
        RECT 962.050 0.010 970.870 4.280 ;
        RECT 971.710 0.010 980.530 4.280 ;
        RECT 981.370 0.010 990.190 4.280 ;
        RECT 991.030 0.010 999.850 4.280 ;
        RECT 1000.690 0.010 1009.510 4.280 ;
        RECT 1010.350 0.010 1019.170 4.280 ;
        RECT 1020.010 0.010 1028.830 4.280 ;
        RECT 1029.670 0.010 1038.490 4.280 ;
        RECT 1039.330 0.010 1048.150 4.280 ;
        RECT 1048.990 0.010 1057.810 4.280 ;
        RECT 1058.650 0.010 1067.470 4.280 ;
        RECT 1068.310 0.010 1077.130 4.280 ;
        RECT 1077.970 0.010 1086.790 4.280 ;
        RECT 1087.630 0.010 1096.450 4.280 ;
        RECT 1097.290 0.010 1106.110 4.280 ;
        RECT 1106.950 0.010 1115.770 4.280 ;
        RECT 1116.610 0.010 1125.430 4.280 ;
        RECT 1126.270 0.010 1135.090 4.280 ;
        RECT 1135.930 0.010 1144.750 4.280 ;
        RECT 1145.590 0.010 1154.410 4.280 ;
        RECT 1155.250 0.010 1164.070 4.280 ;
        RECT 1164.910 0.010 1173.730 4.280 ;
        RECT 1174.570 0.010 1183.390 4.280 ;
        RECT 1184.230 0.010 1193.050 4.280 ;
        RECT 1193.890 0.010 1202.710 4.280 ;
        RECT 1203.550 0.010 1212.370 4.280 ;
        RECT 1213.210 0.010 1222.030 4.280 ;
        RECT 1222.870 0.010 1231.690 4.280 ;
        RECT 1232.530 0.010 1241.350 4.280 ;
        RECT 1242.190 0.010 1251.010 4.280 ;
        RECT 1251.850 0.010 1260.670 4.280 ;
        RECT 1261.510 0.010 1270.330 4.280 ;
        RECT 1271.170 0.010 1279.990 4.280 ;
        RECT 1280.830 0.010 1289.650 4.280 ;
        RECT 1290.490 0.010 1299.310 4.280 ;
        RECT 1300.150 0.010 1308.970 4.280 ;
        RECT 1309.810 0.010 1318.630 4.280 ;
        RECT 1319.470 0.010 1328.290 4.280 ;
        RECT 1329.130 0.010 1337.950 4.280 ;
        RECT 1338.790 0.010 1347.610 4.280 ;
        RECT 1348.450 0.010 1357.270 4.280 ;
        RECT 1358.110 0.010 1366.930 4.280 ;
        RECT 1367.770 0.010 1376.590 4.280 ;
        RECT 1377.430 0.010 1386.250 4.280 ;
        RECT 1387.090 0.010 1395.910 4.280 ;
        RECT 1396.750 0.010 1405.570 4.280 ;
        RECT 1406.410 0.010 1415.230 4.280 ;
        RECT 1416.070 0.010 1424.890 4.280 ;
      LAYER met3 ;
        RECT 10.105 823.480 1371.195 856.625 ;
        RECT 10.105 811.720 1371.195 820.920 ;
        RECT 10.105 773.480 1371.195 809.160 ;
        RECT 10.105 761.720 1371.195 770.920 ;
        RECT 10.105 723.480 1371.195 759.160 ;
        RECT 10.105 711.720 1371.195 720.920 ;
        RECT 10.105 673.480 1371.195 709.160 ;
        RECT 10.105 670.920 324.590 673.480 ;
        RECT 350.200 670.920 674.590 673.480 ;
        RECT 700.200 670.920 1024.590 673.480 ;
        RECT 1050.200 670.920 1371.195 673.480 ;
        RECT 10.105 661.720 1371.195 670.920 ;
        RECT 10.105 623.480 1371.195 659.160 ;
        RECT 10.105 611.720 1371.195 620.920 ;
        RECT 10.105 573.480 1371.195 609.160 ;
        RECT 10.105 561.720 1371.195 570.920 ;
        RECT 10.105 523.480 1371.195 559.160 ;
        RECT 10.105 511.720 1371.195 520.920 ;
        RECT 10.105 473.480 1371.195 509.160 ;
        RECT 10.105 461.720 1371.195 470.920 ;
        RECT 10.105 455.180 1371.195 459.160 ;
        RECT 10.105 423.480 1371.195 452.620 ;
        RECT 10.105 411.720 1371.195 420.920 ;
        RECT 10.105 373.480 1371.195 409.160 ;
        RECT 10.105 361.720 1371.195 370.920 ;
        RECT 10.105 323.480 1371.195 359.160 ;
        RECT 10.105 311.720 1371.195 320.920 ;
        RECT 10.105 273.480 1371.195 309.160 ;
        RECT 10.105 261.720 1371.195 270.920 ;
        RECT 10.105 223.480 1371.195 259.160 ;
        RECT 10.105 211.720 1371.195 220.920 ;
        RECT 10.105 173.480 1371.195 209.160 ;
        RECT 10.105 161.720 1371.195 170.920 ;
        RECT 10.105 123.480 1371.195 159.160 ;
        RECT 10.105 111.720 1371.195 120.920 ;
        RECT 10.105 73.480 1371.195 109.160 ;
        RECT 10.105 61.720 1371.195 70.920 ;
        RECT 10.105 23.480 1371.195 59.160 ;
        RECT 10.105 11.720 1371.195 20.920 ;
        RECT 10.105 0.175 1371.195 9.160 ;
      LAYER met4 ;
        RECT 314.015 0.175 323.110 856.625 ;
        RECT 327.010 0.175 338.110 856.625 ;
        RECT 342.010 0.175 353.110 856.625 ;
        RECT 357.010 0.175 368.110 856.625 ;
        RECT 372.010 0.175 383.110 856.625 ;
        RECT 387.010 0.175 398.110 856.625 ;
        RECT 402.010 0.175 413.110 856.625 ;
        RECT 417.010 0.175 428.110 856.625 ;
        RECT 432.010 0.175 443.110 856.625 ;
        RECT 447.010 0.175 458.110 856.625 ;
        RECT 462.010 0.175 473.110 856.625 ;
        RECT 477.010 0.175 488.110 856.625 ;
        RECT 492.010 0.175 503.110 856.625 ;
        RECT 507.010 0.175 518.110 856.625 ;
        RECT 522.010 0.175 533.110 856.625 ;
        RECT 537.010 0.175 548.110 856.625 ;
        RECT 552.010 0.175 563.110 856.625 ;
        RECT 567.010 0.175 578.110 856.625 ;
        RECT 582.010 0.175 593.110 856.625 ;
        RECT 597.010 0.175 608.110 856.625 ;
        RECT 612.010 0.175 623.110 856.625 ;
        RECT 627.010 0.175 638.110 856.625 ;
        RECT 642.010 0.175 653.110 856.625 ;
        RECT 657.010 0.175 668.110 856.625 ;
        RECT 672.010 0.175 683.110 856.625 ;
        RECT 687.010 0.175 698.110 856.625 ;
        RECT 702.010 0.175 713.110 856.625 ;
        RECT 717.010 0.175 728.110 856.625 ;
        RECT 732.010 0.175 743.110 856.625 ;
        RECT 747.010 0.175 758.110 856.625 ;
        RECT 762.010 0.175 773.110 856.625 ;
        RECT 777.010 0.175 788.110 856.625 ;
        RECT 792.010 0.175 803.110 856.625 ;
        RECT 807.010 0.175 818.110 856.625 ;
        RECT 822.010 0.175 833.110 856.625 ;
        RECT 837.010 0.175 848.110 856.625 ;
        RECT 852.010 0.175 863.110 856.625 ;
        RECT 867.010 0.175 878.110 856.625 ;
        RECT 882.010 0.175 893.110 856.625 ;
        RECT 897.010 0.175 908.110 856.625 ;
        RECT 912.010 0.175 923.110 856.625 ;
        RECT 927.010 0.175 938.110 856.625 ;
        RECT 942.010 0.175 953.110 856.625 ;
        RECT 957.010 0.175 968.110 856.625 ;
        RECT 972.010 0.175 983.110 856.625 ;
        RECT 987.010 0.175 998.110 856.625 ;
        RECT 1002.010 0.175 1013.110 856.625 ;
        RECT 1017.010 0.175 1028.110 856.625 ;
        RECT 1032.010 0.175 1043.110 856.625 ;
        RECT 1047.010 0.175 1058.110 856.625 ;
        RECT 1062.010 0.175 1073.110 856.625 ;
        RECT 1077.010 0.175 1088.110 856.625 ;
        RECT 1092.010 0.175 1103.110 856.625 ;
        RECT 1107.010 0.175 1118.110 856.625 ;
        RECT 1122.010 0.175 1133.110 856.625 ;
        RECT 1137.010 0.175 1148.110 856.625 ;
        RECT 1152.010 0.175 1163.110 856.625 ;
        RECT 1167.010 0.175 1178.110 856.625 ;
        RECT 1182.010 0.175 1193.110 856.625 ;
        RECT 1197.010 0.175 1208.110 856.625 ;
        RECT 1212.010 0.175 1223.110 856.625 ;
        RECT 1227.010 0.175 1238.110 856.625 ;
        RECT 1242.010 0.175 1253.110 856.625 ;
        RECT 1257.010 0.175 1268.110 856.625 ;
        RECT 1272.010 0.175 1283.110 856.625 ;
        RECT 1287.010 0.175 1298.110 856.625 ;
        RECT 1302.010 0.175 1313.110 856.625 ;
        RECT 1317.010 0.175 1328.110 856.625 ;
        RECT 1332.010 0.175 1343.110 856.625 ;
        RECT 1347.010 0.175 1358.110 856.625 ;
        RECT 1362.010 0.175 1365.905 856.625 ;
      LAYER met5 ;
        RECT 872.740 470.100 1352.740 475.100 ;
  END
END CF_SRAM_8192x32
END LIBRARY

